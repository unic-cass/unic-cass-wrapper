magic
tech ihp-sg13g2
magscale 1 2
timestamp 1768335505
<< metal7 >>
rect 70600 372000 84600 386000
rect 91000 372000 105000 386000
rect 111400 372000 125400 386000
rect 131800 372000 145800 386000
rect 152200 372000 166200 386000
rect 172600 372000 186600 386000
rect 193000 372000 207000 386000
rect 213400 372000 227400 386000
rect 233800 372000 247800 386000
rect 254200 372000 268200 386000
rect 274600 372000 288600 386000
rect 295000 372000 309000 386000
rect 315400 372000 329400 386000
rect 14000 315400 28000 329400
rect 372000 315400 386000 329400
rect 14000 295000 28000 309000
rect 372000 295000 386000 309000
rect 14000 274600 28000 288600
rect 372000 274600 386000 288600
rect 14000 254200 28000 268200
rect 372000 254200 386000 268200
rect 14000 233800 28000 247800
rect 372000 233800 386000 247800
rect 14000 213400 28000 227400
rect 372000 213400 386000 227400
rect 14000 193000 28000 207000
rect 372000 193000 386000 207000
rect 14000 172600 28000 186600
rect 372000 172600 386000 186600
rect 14000 152200 28000 166200
rect 372000 152200 386000 166200
rect 14000 131800 28000 145800
rect 372000 131800 386000 145800
rect 14000 111400 28000 125400
rect 372000 111400 386000 125400
rect 14000 91000 28000 105000
rect 372000 91000 386000 105000
rect 14000 70600 28000 84600
rect 372000 70600 386000 84600
rect 70600 14000 84600 28000
rect 91000 14000 105000 28000
rect 111400 14000 125400 28000
rect 131800 14000 145800 28000
rect 152200 14000 166200 28000
rect 172600 14000 186600 28000
rect 193000 14000 207000 28000
rect 213400 14000 227400 28000
rect 233800 14000 247800 28000
rect 254200 14000 268200 28000
rect 274600 14000 288600 28000
rect 295000 14000 309000 28000
rect 315400 14000 329400 28000
use bondpad_70x70  IO_BOND_sg13g2_IOPad_analog_io_0
timestamp 1544794771
transform 1 0 254200 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPad_analog_io_1
timestamp 1544794771
transform 1 0 254200 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPad_io_clock
timestamp 1544794771
transform 1 0 274600 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPad_io_reset
timestamp 1544794771
transform 1 0 274600 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[0\].ui
timestamp 1544794771
transform 0 1 14000 1 0 111400
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[1\].ui
timestamp 1544794771
transform 0 1 14000 1 0 131800
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[2\].ui
timestamp 1544794771
transform 0 1 14000 1 0 152200
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[3\].ui
timestamp 1544794771
transform 0 1 14000 1 0 172600
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[4\].ui
timestamp 1544794771
transform 0 1 14000 1 0 193000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[5\].ui
timestamp 1544794771
transform 0 1 14000 1 0 213400
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[6\].ui
timestamp 1544794771
transform 0 1 14000 1 0 233800
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[7\].ui
timestamp 1544794771
transform 0 1 14000 1 0 254200
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[8\].ui
timestamp 1544794771
transform 0 1 14000 1 0 274600
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[9\].ui
timestamp 1544794771
transform 1 0 111400 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[10\].ui
timestamp 1544794771
transform 1 0 131800 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[11\].ui
timestamp 1544794771
transform 1 0 152200 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[12\].ui
timestamp 1544794771
transform 1 0 172600 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[13\].ui
timestamp 1544794771
transform 1 0 193000 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[14\].ui
timestamp 1544794771
transform 1 0 213400 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[15\].ui
timestamp 1544794771
transform 1 0 233800 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVdd_east
timestamp 1544794771
transform 0 -1 386000 1 0 295000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVdd_north
timestamp 1544794771
transform 1 0 295000 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVdd_south
timestamp 1544794771
transform 1 0 295000 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVdd_west
timestamp 1544794771
transform 0 1 14000 1 0 295000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVss_east
timestamp 1544794771
transform 0 -1 386000 1 0 315400
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVss_north
timestamp 1544794771
transform 1 0 315400 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVss_south
timestamp 1544794771
transform 1 0 315400 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVss_west
timestamp 1544794771
transform 0 1 14000 1 0 315400
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[0\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 111400
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[1\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 131800
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[2\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 152200
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[3\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 172600
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[4\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 193000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[5\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 213400
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[6\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 233800
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[7\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 254200
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[8\].uo
timestamp 1544794771
transform 0 -1 386000 1 0 274600
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[9\].uo
timestamp 1544794771
transform 1 0 111400 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[10\].uo
timestamp 1544794771
transform 1 0 131800 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[11\].uo
timestamp 1544794771
transform 1 0 152200 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[12\].uo
timestamp 1544794771
transform 1 0 172600 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[13\].uo
timestamp 1544794771
transform 1 0 193000 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[14\].uo
timestamp 1544794771
transform 1 0 213400 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[15\].uo
timestamp 1544794771
transform 1 0 233800 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVdd_east
timestamp 1544794771
transform 0 -1 386000 1 0 70600
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVdd_north
timestamp 1544794771
transform 1 0 70600 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVdd_south
timestamp 1544794771
transform 1 0 70600 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVdd_west
timestamp 1544794771
transform 0 1 14000 1 0 70600
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVss_east
timestamp 1544794771
transform 0 -1 386000 1 0 91000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVss_north
timestamp 1544794771
transform 1 0 91000 0 -1 386000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVss_south
timestamp 1544794771
transform 1 0 91000 0 1 14000
box 0 0 14000 14001
use bondpad_70x70  IO_BOND_sg13g2_IOPadVss_west
timestamp 1544794771
transform 0 1 14000 1 0 91000
box 0 0 14000 14001
use sg13g2_Corner  IO_CORNER_NORTH_EAST_INST
timestamp 1716382778
transform -1 0 372000 0 -1 372000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_NORTH_WEST_INST
timestamp 1716382778
transform 1 0 28000 0 -1 372000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_SOUTH_EAST_INST
timestamp 1716382778
transform -1 0 372000 0 1 28000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_SOUTH_WEST_INST
timestamp 1716382778
transform 1 0 28000 0 1 28000
box 1076 1076 36124 36124
use sg13g2_Filler4000  IO_FILL_IO_EAST_0_0
timestamp 1718206866
transform 0 -1 372000 1 0 64000
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_EAST_0_20
timestamp 1718206802
transform 0 -1 372000 1 0 68000
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_0_25
timestamp 1718206786
transform 0 -1 372000 1 0 69000
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_EAST_0_27
timestamp 1716459628
transform 0 -1 372000 1 0 69400
box -100 1076 300 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_1_0
timestamp 1718206866
transform 0 -1 372000 1 0 85600
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_1_20
timestamp 1718206786
transform 0 -1 372000 1 0 89600
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_2_0
timestamp 1718206866
transform 0 -1 372000 1 0 106000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_2_20
timestamp 1718206786
transform 0 -1 372000 1 0 110000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_3_0
timestamp 1718206866
transform 0 -1 372000 1 0 126400
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_3_20
timestamp 1718206786
transform 0 -1 372000 1 0 130400
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_4_0
timestamp 1718206866
transform 0 -1 372000 1 0 146800
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_4_20
timestamp 1718206786
transform 0 -1 372000 1 0 150800
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_5_0
timestamp 1718206866
transform 0 -1 372000 1 0 167200
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_5_20
timestamp 1718206786
transform 0 -1 372000 1 0 171200
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_6_0
timestamp 1718206866
transform 0 -1 372000 1 0 187600
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_6_20
timestamp 1718206786
transform 0 -1 372000 1 0 191600
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_7_0
timestamp 1718206866
transform 0 -1 372000 1 0 208000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_7_20
timestamp 1718206786
transform 0 -1 372000 1 0 212000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_8_0
timestamp 1718206866
transform 0 -1 372000 1 0 228400
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_8_20
timestamp 1718206786
transform 0 -1 372000 1 0 232400
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_9_0
timestamp 1718206866
transform 0 -1 372000 1 0 248800
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_9_20
timestamp 1718206786
transform 0 -1 372000 1 0 252800
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_10_0
timestamp 1718206866
transform 0 -1 372000 1 0 269200
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_10_20
timestamp 1718206786
transform 0 -1 372000 1 0 273200
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_11_0
timestamp 1718206866
transform 0 -1 372000 1 0 289600
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_11_20
timestamp 1718206786
transform 0 -1 372000 1 0 293600
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_12_0
timestamp 1718206866
transform 0 -1 372000 1 0 310000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_12_20
timestamp 1718206786
transform 0 -1 372000 1 0 314000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_EAST_13_0
timestamp 1718206866
transform 0 -1 372000 1 0 330400
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_EAST_13_20
timestamp 1718206802
transform 0 -1 372000 1 0 334400
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_EAST_13_25
timestamp 1718206786
transform 0 -1 372000 1 0 335400
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_EAST_13_27
timestamp 1716459628
transform 0 -1 372000 1 0 335800
box -100 1076 300 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_0_0
timestamp 1718206866
transform 1 0 64000 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_NORTH_0_20
timestamp 1718206802
transform 1 0 68000 0 -1 372000
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_0_25
timestamp 1718206786
transform 1 0 69000 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_NORTH_0_27
timestamp 1716459628
transform 1 0 69400 0 -1 372000
box -100 1076 300 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_1_0
timestamp 1718206866
transform 1 0 85600 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_1_20
timestamp 1718206786
transform 1 0 89600 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_2_0
timestamp 1718206866
transform 1 0 106000 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_2_20
timestamp 1718206786
transform 1 0 110000 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_3_0
timestamp 1718206866
transform 1 0 126400 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_3_20
timestamp 1718206786
transform 1 0 130400 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_4_0
timestamp 1718206866
transform 1 0 146800 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_4_20
timestamp 1718206786
transform 1 0 150800 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_5_0
timestamp 1718206866
transform 1 0 167200 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_5_20
timestamp 1718206786
transform 1 0 171200 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_6_0
timestamp 1718206866
transform 1 0 187600 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_6_20
timestamp 1718206786
transform 1 0 191600 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_7_0
timestamp 1718206866
transform 1 0 208000 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_7_20
timestamp 1718206786
transform 1 0 212000 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_8_0
timestamp 1718206866
transform 1 0 228400 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_8_20
timestamp 1718206786
transform 1 0 232400 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_9_0
timestamp 1718206866
transform 1 0 248800 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_9_20
timestamp 1718206786
transform 1 0 252800 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_10_0
timestamp 1718206866
transform 1 0 269200 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_10_20
timestamp 1718206786
transform 1 0 273200 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_11_0
timestamp 1718206866
transform 1 0 289600 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_11_20
timestamp 1718206786
transform 1 0 293600 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_12_0
timestamp 1718206866
transform 1 0 310000 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_12_20
timestamp 1718206786
transform 1 0 314000 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_NORTH_13_0
timestamp 1718206866
transform 1 0 330400 0 -1 372000
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_NORTH_13_20
timestamp 1718206802
transform 1 0 334400 0 -1 372000
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_NORTH_13_25
timestamp 1718206786
transform 1 0 335400 0 -1 372000
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_NORTH_13_27
timestamp 1716459628
transform 1 0 335800 0 -1 372000
box -100 1076 300 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_0_0
timestamp 1718206866
transform 1 0 64000 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_SOUTH_0_20
timestamp 1718206802
transform 1 0 68000 0 1 28000
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_0_25
timestamp 1718206786
transform 1 0 69000 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_SOUTH_0_27
timestamp 1716459628
transform 1 0 69400 0 1 28000
box -100 1076 300 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_1_0
timestamp 1718206866
transform 1 0 85600 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_1_20
timestamp 1718206786
transform 1 0 89600 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_2_0
timestamp 1718206866
transform 1 0 106000 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_2_20
timestamp 1718206786
transform 1 0 110000 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_3_0
timestamp 1718206866
transform 1 0 126400 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_3_20
timestamp 1718206786
transform 1 0 130400 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_4_0
timestamp 1718206866
transform 1 0 146800 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_4_20
timestamp 1718206786
transform 1 0 150800 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_5_0
timestamp 1718206866
transform 1 0 167200 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_5_20
timestamp 1718206786
transform 1 0 171200 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_6_0
timestamp 1718206866
transform 1 0 187600 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_6_20
timestamp 1718206786
transform 1 0 191600 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_7_0
timestamp 1718206866
transform 1 0 208000 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_7_20
timestamp 1718206786
transform 1 0 212000 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_8_0
timestamp 1718206866
transform 1 0 228400 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_8_20
timestamp 1718206786
transform 1 0 232400 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_9_0
timestamp 1718206866
transform 1 0 248800 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_9_20
timestamp 1718206786
transform 1 0 252800 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_10_0
timestamp 1718206866
transform 1 0 269200 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_10_20
timestamp 1718206786
transform 1 0 273200 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_11_0
timestamp 1718206866
transform 1 0 289600 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_11_20
timestamp 1718206786
transform 1 0 293600 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_12_0
timestamp 1718206866
transform 1 0 310000 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_12_20
timestamp 1718206786
transform 1 0 314000 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_SOUTH_13_0
timestamp 1718206866
transform 1 0 330400 0 1 28000
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_SOUTH_13_20
timestamp 1718206802
transform 1 0 334400 0 1 28000
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_SOUTH_13_25
timestamp 1718206786
transform 1 0 335400 0 1 28000
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_SOUTH_13_27
timestamp 1716459628
transform 1 0 335800 0 1 28000
box -100 1076 300 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_0_0
timestamp 1718206866
transform 0 1 28000 1 0 64000
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_WEST_0_20
timestamp 1718206802
transform 0 1 28000 1 0 68000
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_0_25
timestamp 1718206786
transform 0 1 28000 1 0 69000
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_WEST_0_27
timestamp 1716459628
transform 0 1 28000 1 0 69400
box -100 1076 300 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_1_0
timestamp 1718206866
transform 0 1 28000 1 0 85600
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_1_20
timestamp 1718206786
transform 0 1 28000 1 0 89600
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_2_0
timestamp 1718206866
transform 0 1 28000 1 0 106000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_2_20
timestamp 1718206786
transform 0 1 28000 1 0 110000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_3_0
timestamp 1718206866
transform 0 1 28000 1 0 126400
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_3_20
timestamp 1718206786
transform 0 1 28000 1 0 130400
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_4_0
timestamp 1718206866
transform 0 1 28000 1 0 146800
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_4_20
timestamp 1718206786
transform 0 1 28000 1 0 150800
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_5_0
timestamp 1718206866
transform 0 1 28000 1 0 167200
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_5_20
timestamp 1718206786
transform 0 1 28000 1 0 171200
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_6_0
timestamp 1718206866
transform 0 1 28000 1 0 187600
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_6_20
timestamp 1718206786
transform 0 1 28000 1 0 191600
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_7_0
timestamp 1718206866
transform 0 1 28000 1 0 208000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_7_20
timestamp 1718206786
transform 0 1 28000 1 0 212000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_8_0
timestamp 1718206866
transform 0 1 28000 1 0 228400
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_8_20
timestamp 1718206786
transform 0 1 28000 1 0 232400
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_9_0
timestamp 1718206866
transform 0 1 28000 1 0 248800
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_9_20
timestamp 1718206786
transform 0 1 28000 1 0 252800
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_10_0
timestamp 1718206866
transform 0 1 28000 1 0 269200
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_10_20
timestamp 1718206786
transform 0 1 28000 1 0 273200
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_11_0
timestamp 1718206866
transform 0 1 28000 1 0 289600
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_11_20
timestamp 1718206786
transform 0 1 28000 1 0 293600
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_12_0
timestamp 1718206866
transform 0 1 28000 1 0 310000
box -124 1076 4124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_12_20
timestamp 1718206786
transform 0 1 28000 1 0 314000
box -124 1076 524 35600
use sg13g2_Filler4000  IO_FILL_IO_WEST_13_0
timestamp 1718206866
transform 0 1 28000 1 0 330400
box -124 1076 4124 35600
use sg13g2_Filler1000  IO_FILL_IO_WEST_13_20
timestamp 1718206802
transform 0 1 28000 1 0 334400
box -124 1076 1124 35600
use sg13g2_Filler400  IO_FILL_IO_WEST_13_25
timestamp 1718206786
transform 0 1 28000 1 0 335400
box -124 1076 524 35600
use sg13g2_Filler200  IO_FILL_IO_WEST_13_27
timestamp 1716459628
transform 0 1 28000 1 0 335800
box -100 1076 300 35600
use sg13g2_IOPadAnalog  sg13g2_IOPad_analog_io_0
timestamp 1718205910
transform 1 0 253200 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadAnalog  sg13g2_IOPad_analog_io_1
timestamp 1718205910
transform 1 0 253200 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPad_io_clock
timestamp 1716382777
transform 1 0 273600 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPad_io_reset
timestamp 1716382777
transform 1 0 273600 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[0\].ui
timestamp 1716382777
transform 0 1 28000 1 0 110400
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[1\].ui
timestamp 1716382777
transform 0 1 28000 1 0 130800
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[2\].ui
timestamp 1716382777
transform 0 1 28000 1 0 151200
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[3\].ui
timestamp 1716382777
transform 0 1 28000 1 0 171600
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[4\].ui
timestamp 1716382777
transform 0 1 28000 1 0 192000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[5\].ui
timestamp 1716382777
transform 0 1 28000 1 0 212400
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[6\].ui
timestamp 1716382777
transform 0 1 28000 1 0 232800
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[7\].ui
timestamp 1716382777
transform 0 1 28000 1 0 253200
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[8\].ui
timestamp 1716382777
transform 0 1 28000 1 0 273600
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[9\].ui
timestamp 1716382777
transform 1 0 110400 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[10\].ui
timestamp 1716382777
transform 1 0 130800 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[11\].ui
timestamp 1716382777
transform 1 0 151200 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[12\].ui
timestamp 1716382777
transform 1 0 171600 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[13\].ui
timestamp 1716382777
transform 1 0 192000 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[14\].ui
timestamp 1716382777
transform 1 0 212400 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[15\].ui
timestamp 1716382777
transform 1 0 232800 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIOVdd  sg13g2_IOPadIOVdd_east
timestamp 1716382778
transform 0 -1 372000 1 0 294000
box -124 0 16124 35600
use sg13g2_IOPadIOVdd  sg13g2_IOPadIOVdd_north
timestamp 1716382778
transform 1 0 294000 0 -1 372000
box -124 0 16124 35600
use sg13g2_IOPadIOVdd  sg13g2_IOPadIOVdd_south
timestamp 1716382778
transform 1 0 294000 0 1 28000
box -124 0 16124 35600
use sg13g2_IOPadIOVdd  sg13g2_IOPadIOVdd_west
timestamp 1716382778
transform 0 1 28000 1 0 294000
box -124 0 16124 35600
use sg13g2_IOPadIOVss  sg13g2_IOPadIOVss_east
timestamp 1716382777
transform 0 -1 372000 1 0 314400
box -124 0 16124 35600
use sg13g2_IOPadIOVss  sg13g2_IOPadIOVss_north
timestamp 1716382777
transform 1 0 314400 0 -1 372000
box -124 0 16124 35600
use sg13g2_IOPadIOVss  sg13g2_IOPadIOVss_south
timestamp 1716382777
transform 1 0 314400 0 1 28000
box -124 0 16124 35600
use sg13g2_IOPadIOVss  sg13g2_IOPadIOVss_west
timestamp 1716382777
transform 0 1 28000 1 0 314400
box -124 0 16124 35600
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[0\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 110400
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[1\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 130800
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[2\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 151200
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[3\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 171600
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[4\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 192000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[5\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 212400
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[6\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 232800
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[7\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 253200
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[8\].uo
timestamp 1716382777
transform 0 -1 372000 1 0 273600
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[9\].uo
timestamp 1716382777
transform 1 0 110400 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[10\].uo
timestamp 1716382777
transform 1 0 130800 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[11\].uo
timestamp 1716382777
transform 1 0 151200 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[12\].uo
timestamp 1716382777
transform 1 0 171600 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[13\].uo
timestamp 1716382777
transform 1 0 192000 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[14\].uo
timestamp 1716382777
transform 1 0 212400 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[15\].uo
timestamp 1716382777
transform 1 0 232800 0 -1 372000
box -124 0 16124 36000
use sg13g2_IOPadVdd  sg13g2_IOPadVdd_east
timestamp 1716382777
transform 0 -1 372000 1 0 69600
box -124 0 16124 35600
use sg13g2_IOPadIOVdd  sg13g2_IOPadVdd_north
timestamp 1716382778
transform 1 0 69600 0 -1 372000
box -124 0 16124 35600
use sg13g2_IOPadVdd  sg13g2_IOPadVdd_south
timestamp 1716382777
transform 1 0 69600 0 1 28000
box -124 0 16124 35600
use sg13g2_IOPadVdd  sg13g2_IOPadVdd_west
timestamp 1716382777
transform 0 1 28000 1 0 69600
box -124 0 16124 35600
use sg13g2_IOPadVss  sg13g2_IOPadVss_east
timestamp 1716382777
transform 0 -1 372000 1 0 90000
box -124 0 16124 35600
use sg13g2_IOPadIOVss  sg13g2_IOPadVss_north
timestamp 1716382777
transform 1 0 90000 0 -1 372000
box -124 0 16124 35600
use sg13g2_IOPadVss  sg13g2_IOPadVss_south
timestamp 1716382777
transform 1 0 90000 0 1 28000
box -124 0 16124 35600
use sg13g2_IOPadVss  sg13g2_IOPadVss_west
timestamp 1716382777
transform 0 1 28000 1 0 90000
box -124 0 16124 35600
<< labels >>
flabel metal7 s 14000 295000 28000 309000 0 FreeSans 102400 0 0 0 IOVDD
port 0 nsew power input
flabel metal7 s 295000 372000 309000 386000 0 FreeSans 102400 0 0 0 IOVDD
port 1 nsew power input
flabel metal7 s 70600 372000 84600 386000 0 FreeSans 102400 0 0 0 IOVDD
port 2 nsew power input
flabel metal7 s 372000 295000 386000 309000 0 FreeSans 102400 0 0 0 IOVDD
port 3 nsew power input
flabel metal7 s 295000 14000 309000 28000 0 FreeSans 102400 0 0 0 IOVDD
port 4 nsew power input
flabel metal7 s 14000 315400 28000 329400 0 FreeSans 102400 0 0 0 IOVSS
port 5 nsew ground input
flabel metal7 s 315400 372000 329400 386000 0 FreeSans 102400 0 0 0 IOVSS
port 6 nsew ground input
flabel metal7 s 91000 372000 105000 386000 0 FreeSans 102400 0 0 0 IOVSS
port 7 nsew ground input
flabel metal7 s 372000 315400 386000 329400 0 FreeSans 102400 0 0 0 IOVSS
port 8 nsew ground input
flabel metal7 s 315400 14000 329400 28000 0 FreeSans 102400 0 0 0 IOVSS
port 9 nsew ground input
flabel metal7 s 14000 70600 28000 84600 0 FreeSans 102400 0 0 0 VDD
port 10 nsew power input
flabel metal7 s 372000 70600 386000 84600 0 FreeSans 102400 0 0 0 VDD
port 11 nsew power input
flabel metal7 s 70600 14000 84600 28000 0 FreeSans 102400 0 0 0 VDD
port 12 nsew power input
flabel metal7 s 14000 91000 28000 105000 0 FreeSans 102400 0 0 0 VSS
port 13 nsew ground input
flabel metal7 s 372000 91000 386000 105000 0 FreeSans 102400 0 0 0 VSS
port 14 nsew ground input
flabel metal7 s 91000 14000 105000 28000 0 FreeSans 102400 0 0 0 VSS
port 15 nsew ground input
flabel metal7 s 254200 14000 268200 28000 0 FreeSans 102400 0 0 0 analog_io_0
port 16 nsew signal bidirectional
flabel metal7 s 254200 372000 268200 386000 0 FreeSans 102400 0 0 0 analog_io_1
port 17 nsew signal bidirectional
flabel metal7 s 274600 14000 288600 28000 0 FreeSans 102400 0 0 0 io_clock_PAD
port 18 nsew signal bidirectional
flabel metal7 s 274600 372000 288600 386000 0 FreeSans 102400 0 0 0 io_reset_PAD
port 19 nsew signal bidirectional
flabel metal7 s 14000 111400 28000 125400 0 FreeSans 102400 0 0 0 ui_PAD[0]
port 20 nsew signal bidirectional
flabel metal7 s 131800 14000 145800 28000 0 FreeSans 102400 0 0 0 ui_PAD[10]
port 21 nsew signal bidirectional
flabel metal7 s 152200 14000 166200 28000 0 FreeSans 102400 0 0 0 ui_PAD[11]
port 22 nsew signal bidirectional
flabel metal7 s 172600 14000 186600 28000 0 FreeSans 102400 0 0 0 ui_PAD[12]
port 23 nsew signal bidirectional
flabel metal7 s 193000 14000 207000 28000 0 FreeSans 102400 0 0 0 ui_PAD[13]
port 24 nsew signal bidirectional
flabel metal7 s 213400 14000 227400 28000 0 FreeSans 102400 0 0 0 ui_PAD[14]
port 25 nsew signal bidirectional
flabel metal7 s 233800 14000 247800 28000 0 FreeSans 102400 0 0 0 ui_PAD[15]
port 26 nsew signal bidirectional
flabel metal7 s 14000 131800 28000 145800 0 FreeSans 102400 0 0 0 ui_PAD[1]
port 27 nsew signal bidirectional
flabel metal7 s 14000 152200 28000 166200 0 FreeSans 102400 0 0 0 ui_PAD[2]
port 28 nsew signal bidirectional
flabel metal7 s 14000 172600 28000 186600 0 FreeSans 102400 0 0 0 ui_PAD[3]
port 29 nsew signal bidirectional
flabel metal7 s 14000 193000 28000 207000 0 FreeSans 102400 0 0 0 ui_PAD[4]
port 30 nsew signal bidirectional
flabel metal7 s 14000 213400 28000 227400 0 FreeSans 102400 0 0 0 ui_PAD[5]
port 31 nsew signal bidirectional
flabel metal7 s 14000 233800 28000 247800 0 FreeSans 102400 0 0 0 ui_PAD[6]
port 32 nsew signal bidirectional
flabel metal7 s 14000 254200 28000 268200 0 FreeSans 102400 0 0 0 ui_PAD[7]
port 33 nsew signal bidirectional
flabel metal7 s 14000 274600 28000 288600 0 FreeSans 102400 0 0 0 ui_PAD[8]
port 34 nsew signal bidirectional
flabel metal7 s 111400 14000 125400 28000 0 FreeSans 102400 0 0 0 ui_PAD[9]
port 35 nsew signal bidirectional
flabel metal7 s 372000 111400 386000 125400 0 FreeSans 102400 0 0 0 uo_PAD[0]
port 36 nsew signal bidirectional
flabel metal7 s 131800 372000 145800 386000 0 FreeSans 102400 0 0 0 uo_PAD[10]
port 37 nsew signal bidirectional
flabel metal7 s 152200 372000 166200 386000 0 FreeSans 102400 0 0 0 uo_PAD[11]
port 38 nsew signal bidirectional
flabel metal7 s 172600 372000 186600 386000 0 FreeSans 102400 0 0 0 uo_PAD[12]
port 39 nsew signal bidirectional
flabel metal7 s 193000 372000 207000 386000 0 FreeSans 102400 0 0 0 uo_PAD[13]
port 40 nsew signal bidirectional
flabel metal7 s 213400 372000 227400 386000 0 FreeSans 102400 0 0 0 uo_PAD[14]
port 41 nsew signal bidirectional
flabel metal7 s 233800 372000 247800 386000 0 FreeSans 102400 0 0 0 uo_PAD[15]
port 42 nsew signal bidirectional
flabel metal7 s 372000 131800 386000 145800 0 FreeSans 102400 0 0 0 uo_PAD[1]
port 43 nsew signal bidirectional
flabel metal7 s 372000 152200 386000 166200 0 FreeSans 102400 0 0 0 uo_PAD[2]
port 44 nsew signal bidirectional
flabel metal7 s 372000 172600 386000 186600 0 FreeSans 102400 0 0 0 uo_PAD[3]
port 45 nsew signal bidirectional
flabel metal7 s 372000 193000 386000 207000 0 FreeSans 102400 0 0 0 uo_PAD[4]
port 46 nsew signal bidirectional
flabel metal7 s 372000 213400 386000 227400 0 FreeSans 102400 0 0 0 uo_PAD[5]
port 47 nsew signal bidirectional
flabel metal7 s 372000 233800 386000 247800 0 FreeSans 102400 0 0 0 uo_PAD[6]
port 48 nsew signal bidirectional
flabel metal7 s 372000 254200 386000 268200 0 FreeSans 102400 0 0 0 uo_PAD[7]
port 49 nsew signal bidirectional
flabel metal7 s 372000 274600 386000 288600 0 FreeSans 102400 0 0 0 uo_PAD[8]
port 50 nsew signal bidirectional
flabel metal7 s 111400 372000 125400 386000 0 FreeSans 102400 0 0 0 uo_PAD[9]
port 51 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 400000 400000
<< end >>
